

package seq_pkg;
   import uvm_pkg::*;
`include "uvm_macros.svh"
`include "riscv_seq_item.svh"
`include "riscv_seqr.sv"
`include "sequence_base.svh"

endpackage
